open corebase
open coreext
open layers
open tensorm
open corecuda
open rangem

type graph_body = tensor d3 cem.prob * cem.model * cem.trace_state

inl trace_and_play_ forall inp out.
        (is_train : bool) // The sampling behavior differs depending on whether the training is being done.
        rng
        (model : model graph_body)
        (sizes : cem.sizes)
        (exists mid. input : exists mid. (inp -> mid) * pickler.pu mid) 
        (output : int -> out) 
        ~({player_id}, data : {player_id : cem.player_id} * inp) =
    // Get the ensemble,block and thread dimensions based on the output tensor.
    inl ensemble,block,thread,inner = (key_extract model .output_probs : tensor d4 float).dim
    inl () = // Assert that all the dimensions are right.
        assert (block = blocks_per_grid()) "The second dimension of the output tensor has to equal the number of blocks per grid."
        assert (thread = threads_per_block()) "The third dimension of the output tensor has to equal number threads per block."
        inl block',thread',_ = (key_extract model .input : tensor d3 float).dim
        assert ((block,thread) = (block',thread')) "The first two dimensions of the input tensor have to match number of blocks per grid and number of threads per block respectively."

    // Extract the input tensor.
    inl x = (key_extract model .input : tensor d3 float)
    assert (block = fst x.dim) "The first dimension of the input tensor has to equal the number of blocks per grid."
    inl x = x |> apply block_index()
    assert (thread = fst x.dim) "The second dimension of the input tensor has to equal number threads per block."

    // Sets the input tensor to 0.
    loop.projective threads_in_block(x.dim) fun i =>
        tensor_set i 0 x

    __syncthreads()

    // Serializes the data into the input tensor.
    inl () =
        open pickler
        inl tns_input = apply thread_index() x
        snd input .pickle (fst input data) (0,tns_input |> ptr_at_current_offset)

    __syncthreads()

    // Creates the layer state.
    inl ls = create_layer_state rng

    // Runs the model on the inputs.
    loop.linear ensemble fun ensemble =>
        graph_run_device model ls {ensemble}

    __syncthreads()

    // Extract the cem model.
    inl cem_model = (key_extract model .cem_model : cem.model)

    // Extract the output index and the sampling probability for it.
    inl sampling,action_id =
        inl ensemble_id : int = 
            if is_train then
                // The ensemble id is held steady between the `apply_updates` calls.
                tensor_index {} cem_model.exploratory_ensemble_id
            else
                // Generates a random ensemble_id and shares it across all the threads in the block.
                random.int_range {from=0; nearTo=sizes.ensemble_id} rng
                |> transposing_loop.shuffle 0

        cem.get_action rng model ensemble_id
        // Shares the action_id across all the threads in the block.
        |> transposing_loop.shuffle 0

    // Extract the cem trace state model.
    inl cem_trace_state = (key_extract model .cem_trace_state : cem.trace_state)
    
    // Index of the thread in the grid.
    inl thread_id = rangem.threads_in_grid().from

    loop.linear ensemble fun ensemble_id =>
        // Calculate the policy probability for the given action.
        inl policy = cem.get_policy_probs model ensemble_id action_id
        cem.update_trace_state_path_probs cem_trace_state {thread_id ensemble_id player_id} ({policy sampling}, action_id)

    output action_id

inl run_ forall inp out.
        rng
        (model : model graph_body)
        (exists mid. input : exists mid. (inp -> mid) * pickler.pu mid)
        (output : int -> out)
        ~(data : inp) =
    // Get the ensemble,block and thread dimensions based on the output tensor.
    inl ensemble,block,thread,inner = (key_extract model .output_probs : tensor d4 float).dim
    inl () = // Assert that all the dimensions are right.
        assert (block = blocks_per_grid()) "The second dimension of the output tensor has to equal the number of blocks per grid."
        assert (thread = threads_per_block()) "The third dimension of the output tensor has to equal number threads per block."
        inl block',thread',_ = (key_extract model .input : tensor d3 float).dim
        assert ((block,thread) = (block',thread')) "The first two dimensions of the input tensor have to match number of blocks per grid and number of threads per block respectively."

    // Extract the input tensor.
    inl x = (key_extract model .input : tensor d3 float)
    assert (block = fst x.dim) "The first dimension of the input tensor has to equal the number of blocks per grid."
    inl x = x |> apply block_index()
    assert (thread = fst x.dim) "The second dimension of the input tensor has to equal number threads per block."

    // Sets the input tensor to 0.
    loop.projective threads_in_block(x.dim) fun i =>
        tensor_set i 0 x

    __syncthreads()

    // Serializes the data into the input tensor.
    inl () =
        open pickler
        inl tns_input = apply thread_index() x
        snd input .pickle (fst input data) (0,tns_input |> ptr_at_current_offset)

    __syncthreads()

    // TODO: Might have to change this to a loop once we do RNNs.

    // Randomly pick an ensemble id for each thread.
    inl ensemble_id : int = 
        random.int_range {from=0; nearTo=ensemble} rng
        |> transposing_loop.shuffle 0

    // Creates the layer state.
    inl ls = create_layer_state rng

    // Runs the model on the inputs.
    graph_run_device model ls {ensemble=ensemble_id}

    __syncthreads()
    
    output (cem.get_action rng model ensemble_id |> snd)

nominal cem_game_graph inp out =
    {
        graph : graph graph_body
        sizes : cem.sizes
        input : exists t. (inp -> t) * pickler.pu t
        output : int -> out
    }

nominal cem_game_model inp out = 
    {
        model : model graph_body
        sizes : cem.sizes
        input : exists t. (inp -> t) * pickler.pu t
        output : int -> out
    }

inl run forall inp out. rng (cem_game_model {model input output} : cem_game_model inp out) = run_ rng model input output

inl to_model_ptrs forall a b. (cem_game_model {model} : cem_game_model a b) : layers.model_ptrs .cem = model_to_model_ptrs model
inl from_model_ptrs forall inp out. 
        (cem_game_graph {graph sizes input output} : cem_game_graph inp out) 
        (x : layers.model_ptrs .cem)
        : cem_game_model inp out = 
    inl model = model_ptrs_to_model graph x
    cem_game_model { model sizes input output }

inl init forall a b. (cem_game_graph {graph sizes input output} : cem_game_graph a b) : cem_game_model a b = 
    inl model = create_model graph
    pass_init model
    cem_game_model { input sizes output model }

// Applies the index of the thread in the grid.
inl extract_log_path_probs forall inp out. 
        (cem_game_model {model sizes} : cem_game_model inp out) 
        : tensor (path_probs.ensemble_id * path_probs.player_id) path_probs.log_path_prob =
    (key_extract model .cem_trace_state : cem.trace_state).log_path_probs
    |> reorder (fun ensemble_id,thread_id,player_id => thread_id,ensemble_id,player_id)
    |> apply rangem.threads_in_grid().from

inl trace_and_train forall inp out. rng (cem_game_model {model sizes input output} : cem_game_model inp out) = 
    trace_and_play_ true rng model sizes input output

inl trace_and_play forall inp out. rng (cem_game_model {model sizes input output} : cem_game_model inp out) = 
    trace_and_play_ false rng model sizes input output

// Calculates the policy and the value array updates.
// Also resets the trace state afterwards.
inl calculate_updates forall dim a b.
        (cem_game_model {model sizes} : _ a b)
        (reward : sa dim cem.reward) =
    // Since we aren't using the output_world_id we'll pass `ensemble=0` instead of extracting the other nodes one by one.
    inl _, cem_model, trace_state : graph_body = layers.graph_extract model {ensemble=0 : int}
    cem.calculate_updates cem_model trace_state reward

// Resets the trace state.
inl reset_trace_state forall a b. (cem_game_model {model sizes} : _ a b) =
    inl trace_state = (key_extract model .cem_trace_state : cem.trace_state)
    cem.reset_trace_state trace_state

// Applies the policy and the value array updates.
// Clamps the average policy vector if applicable.
// Also randomizes the `exploratory_ensemble_id`.
inl apply_updates forall a b. grid rng (cem_game_model {model} : _ a b) =
    inl x : list (cem_weight_layer_dual float) = key_extract_list model .cem_weight_layer_dual
    inl l : list cem.weights = x |> listm.map (fun a,b => exists a,b)
    inl _, cem_model, trace_state : graph_body = layers.graph_extract model {ensemble=0 : int}
    cem.apply_updates rng grid l cem_model