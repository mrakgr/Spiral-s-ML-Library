open corebase
open coreext
open layers
open tensorm
open corecuda
open rangem

inl print0 msg =
    if rangem.threads_in_grid().from = 0 then
        console.write_ln msg
    __syncwarp()

type graph_body = tensor d2 uint * cfr.model * cfr.trace * cfr.trace_state

inl trace_and_play_ forall inp out.
        (is_train : bool) // The sampling behavior differs depending on whether the training is being done.
        rng
        (model : model graph_body)
        (sizes : cfr.sizes)
        (action_mask : primitives.row_config -> f32 -> i32 -> i32 -> bool)
        (exists mid. input : exists mid. (inp -> mid) * pickler.pu mid) 
        (output : int -> out) 
        ~({player_id}, data : {player_id : cfr.player_id} * inp) =

    // Get the ensemble,block and thread dimensions based on the output tensor.
    inl ensemble,block,thread = (key_extract model .output_world_id : tensor d3 uint).dim
    inl () = // Assert that all the dimensions are right.
        assert (block = blocks_per_grid()) "The second dimension of the output tensor has to equal the number of blocks per grid."
        assert (thread = threads_per_block()) "The third dimension of the output tensor has to equal number threads per block."
        inl block',thread',_ = (key_extract model .input : tensor d3 float).dim
        assert ((block,thread) = (block',thread')) "The first two dimensions of the input tensor have to match number of blocks per grid and number of threads per block respectively."

    // Extract the input tensor.
    inl x = (key_extract model .input : tensor d3 float)
    assert (block = fst x.dim) "The first dimension of the input tensor has to equal the number of blocks per grid."
    inl x = x |> apply block_index()
    assert (thread = fst x.dim) "The second dimension of the input tensor has to equal number threads per block."


    // Sets the input tensor to 0.
    loop.projective threads_in_block(x.dim) fun i =>
        tensor_set i 0 x

    barrier_cta_sync 0

    // Serializes the data into the input tensor.
    inl () =
        open pickler
        inl tns_input = apply thread_index() x
        snd input .pickle (fst input data) (0,tns_input |> ptr_at_current_offset)

    barrier_cta_sync 0

    // Creates the layer state.
    inl ls = create_layer_state rng

    // Runs the model on the inputs.
    loop.linear ensemble fun ensemble =>
        graph_run_device model ls {ensemble}

    barrier_cta_sync 0

    // Extract the CFR model.
    inl cfr_model = (key_extract model .cfr_model : cfr.model)

    // Extract the output index and the sampling probability for it.
    inl sampling,action_id = 
        inl ensemble_id : int = 
            if is_train then
                // The ensemble id is held steady between the `apply_updates` calls.
                tensor_index {} cfr_model.exploratory_ensemble_id
            else
                // Generates a random ensemble_id and shares it across all the threads in the block.
                random.int_range {from=0; nearTo=sizes.ensemble_id} rng
                |> transposing_loop.shuffle 0

        // Extract the hash of the input state for the CFR model.
        inl world_id =
            (key_extract model .output_world_id : tensor d3 uint)
            |> tensor_index (ensemble_id, block_index(), thread_index())

        cfr.get_action rng action_mask cfr_model (ensemble_id, conv world_id)
        // Shares the action_id across all the threads in the block.
        |> transposing_loop.shuffle 0

    // Extract the CFR trace state model.
    inl cfr_trace_state = (key_extract model .cfr_trace_state : cfr.trace_state)
    
    // Extract the CFR trace.
    inl cfr_trace = (key_extract model .cfr_trace : cfr.trace)

    // Index of the thread in the grid.
    inl thread_id = rangem.threads_in_grid().from

    loop.linear ensemble fun ensemble_id =>
        // Extract the hash of the input state for the CFR model.
        inl world_id =
            (key_extract model .output_world_id : tensor d3 uint)
            |> tensor_index (ensemble_id, block_index(), thread_index())
            |> conv


        // Calculate the policy probability for the given action.
        inl policy = 
            if is_train then
                // During training the policy is the current policy.
                cfr.get_policy_probs action_mask cfr_model (ensemble_id, world_id) action_id
            else
                // During evaluation the policy is the average policy.
                cfr.get_average_probs action_mask cfr_model (ensemble_id, world_id) action_id

        if is_train then
            // Pushes the data into the trace.
            cfr.push_trace cfr_trace cfr_trace_state {thread_id ensemble_id world_id player_id} ({policy sampling}, action_id)
        else
            // During eval it only updates the path probabilities for the state. It does not push data into the trace to save computation.
            cfr.update_trace_state_path_probs cfr_trace_state {thread_id ensemble_id player_id} ({policy sampling}, action_id)

    output action_id

inl run_ forall inp out.
        rng
        (model : model graph_body)
        (action_mask : primitives.row_config -> f32 -> i32 -> i32 -> bool)
        (exists mid. input : exists mid. (inp -> mid) * pickler.pu mid) 
        (output : int -> out) 
        (data : inp) =

    // Get the ensemble,block and thread dimensions based on the output tensor.
    inl ensemble,block,thread = (key_extract model .output_world_id : tensor d3 uint).dim
    inl () = // Assert that all the dimensions are right.
        assert (block = blocks_per_grid()) "The second dimension of the output tensor has to equal the number of blocks per grid."
        assert (thread = threads_per_block()) "The third dimension of the output tensor has to equal number threads per block."
        inl block',thread',_ = (key_extract model .input : tensor d3 float).dim
        assert ((block,thread) = (block',thread')) "The first two dimensions of the input tensor have to match number of blocks per grid and number of threads per block respectively."

    // Extract the input tensor.
    inl x = (key_extract model .input : tensor d3 float)
    assert (block = fst x.dim) "The first dimension of the input tensor has to equal the number of blocks per grid."
    inl x = x |> apply block_index()
    assert (thread = fst x.dim) "The second dimension of the input tensor has to equal number threads per block."

    // Sets the input tensor to 0.
    loop.projective threads_in_block(x.dim) fun i =>
        tensor_set i 0 x

    barrier_cta_sync 0

    // Serializes the data into the input tensor.
    inl () =
        open pickler
        inl tns_input = apply thread_index() x
        snd input .pickle (fst input data) (0,tns_input |> ptr_at_current_offset)

    barrier_cta_sync 0

    // Randomly pick an ensemble id for each thread.
    inl ensemble_id : int = 
        random.int_range {from=0; nearTo=ensemble} ls.rng
        |> transposing_loop.shuffle 0

    // Creates the layer state.
    inl ls = create_layer_state rng

    // Runs the model on the inputs.
    graph_run_device model ls {ensemble=ensemble_id}

    barrier_cta_sync 0

    // Extract the hash of the input state.
    inl world_id =
        (key_extract model .output_world_id : tensor d3 uint)
        |> tensor_index (ensemble_id, block_index(), thread_index())

    // Extract the CFR model.
    inl cfr_model = (key_extract model .cfr_model : cfr.model)

    // Extract the output index.
    inl _,output_id = cfr.get_action rng action_mask cfr_model (ensemble_id, conv world_id)

    output output_id

nominal cfr_game_graph inp out =
    {
        graph : graph graph_body
        sizes : cfr.sizes
        action_mask : primitives.row_config -> f32 -> i32 -> i32 -> bool
        input : exists t. (inp -> t) * pickler.pu t
        output : int -> out
    }

nominal cfr_game_model inp out = 
    {
        model : model graph_body
        sizes : cfr.sizes
        action_mask : primitives.row_config -> f32 -> i32 -> i32 -> bool
        input : exists t. (inp -> t) * pickler.pu t
        output : int -> out
    }

// Integrates all the path probabilities. Integrates out the ensemble id before multiplyting the player probabilities.
// 
// Pseudo-code: 
// prod (fun player_id => sum (fun ensemble_id => p(player_id,ensemble_id)))
inl extract_integrated_path_prob forall inp out. (cfr_game_model {model sizes} : cfr_game_model inp out) : cfr.prob =
    inl log_path_probs = 
        (key_extract model .cfr_trace_state : cfr.trace_state).log_path_probs
        |> reorder (fun ensemble_id,thread_id,player_id => thread_id,player_id,ensemble_id)
        |> apply rangem.threads_in_grid().from
    loop.for {from=0; nearTo=sizes.player_id} (fun player_id s =>
        inl log_path_probs = apply player_id log_path_probs
        s * loop.for {from=0; nearTo=sizes.ensemble_id} (fun ensemble_id s => 
            inl {policy sampling} = tensor_index ensemble_id log_path_probs
            s + exp (policy - sampling)
            ) 0
        ) 1
    |> conv

// Excludes the ensemble from the path probability calculations.
inl extract_integrated_path_prob_excluding forall inp out. (cfr_game_model {model sizes} : cfr_game_model inp out) {ensemble_id} : cfr.prob =
    inl log_path_probs = 
        (key_extract model .cfr_trace_state : cfr.trace_state).log_path_probs
        |> reorder (fun ensemble_id,thread_id,player_id => thread_id,player_id,ensemble_id)
        |> apply rangem.threads_in_grid().from
    loop.for {from=0; nearTo=sizes.player_id} (fun player_id s =>
        inl log_path_probs = apply player_id log_path_probs
        s * loop.for {from=0; nearTo=sizes.ensemble_id} (fun ensemble_id' s => 
            inl {policy sampling} = tensor_index ensemble_id' log_path_probs
            inl p = exp (policy - sampling)
            s + (if ensemble_id <> ensemble_id' then p else 0)
            ) 0
        ) 1
    |> conv

// Extracts the path probability conditioned on an ensemble_id.
inl extract_ensemble_path_prob forall inp out. (m : cfr_game_model inp out) ensemble_id =
    extract_integrated_path_prob m - extract_integrated_path_prob_excluding m ensemble_id

inl run forall inp out. rng (cfr_game_model {model action_mask input output} : cfr_game_model inp out) = run_ rng model action_mask input output
inl trace_and_train forall inp out. rng (cfr_game_model {model sizes action_mask input output} : cfr_game_model inp out) = 
    trace_and_play_ true rng model sizes action_mask input output

inl trace_and_play forall inp out. rng (cfr_game_model {model sizes action_mask input output} : cfr_game_model inp out) = 
    trace_and_play_ false rng model sizes action_mask input output

inl to_model_data forall a b. (cfr_game_model {model} : cfr_game_model a b) : layers.model_data = model_to_model_data model
inl from_model_data forall inp out.
        (cfr_game_graph {graph sizes input output action_mask} : cfr_game_graph inp out) 
        (x : layers.model_data) 
        : cfr_game_model inp out = 
    inl model = model_data_to_model graph x
    cfr_game_model {model sizes action_mask input output}

inl init forall a b. (cfr_game_graph {graph sizes action_mask input output} : cfr_game_graph a b) : cfr_game_model a b = 
    inl model = create_model graph
    param_init model
    cfr_game_model { sizes input output action_mask model }

// Calculates the policy and the value array updates.
// Also resets the trace state afterwards.
inl calculate_updates forall dim a b.
        (cfr_game_model {model sizes action_mask} : _ a b)
        (reward : sa dim cfr.reward) =
    // Since we aren't using the output_world_id we'll pass `ensemble=0` instead of extracting the other nodes one by one.
    inl _, cfr_model, trace, trace_state : graph_body = layers.graph_extract model {ensemble=0 : int}
    loop.linear sizes.ensemble_id fun ensemble_id =>
        cfr.calculate_updates action_mask sizes cfr_model trace trace_state ensemble_id reward

// Resets the trace state.
inl reset_trace_state forall a b. (cfr_game_model {model sizes} : _ a b) =
    inl trace_state = (key_extract model .cfr_trace_state : cfr.trace_state)
    loop.linear sizes.ensemble_id fun ensemble_id =>
        cfr.reset_trace_state trace_state ensemble_id

// Applies the policy and the value array updates.
// Clamps the average policy vector if applicable.
// Also randomizes the `exploratory_ensemble_id`.
inl apply_updates forall a b. grid rng (cfr_game_model {model} : _ a b) =
    inl _, cfr_model, trace, trace_state : graph_body = layers.graph_extract model {ensemble=0 : int}
    cfr.apply_updates grid rng cfr_model